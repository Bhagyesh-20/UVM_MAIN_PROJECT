0 | rst_n=0 | Addr=0000 | cmd_n=1 | RDnWR=0 | DataIn=00000000 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=0 | RA=0 | CA=0 | cs_n=0
#                   20 | rst_n=1 | Addr=0000 | cmd_n=1 | RDnWR=0 | DataIn=00000000 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=0 | RA=0 | CA=0 | cs_n=0
#                   25 | rst_n=1 | Addr=0000 | cmd_n=1 | RDnWR=0 | DataIn=00000000 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=4 | DataOutVld=1 | RA=0 | CA=0 | cs_n=0
#                   35 | rst_n=1 | Addr=0000 | cmd_n=1 | RDnWR=0 | DataIn=00000000 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=1 | RA=0 | CA=0 | cs_n=0
#                   45 | rst_n=1 | Addr=0000 | cmd_n=1 | RDnWR=0 | DataIn=00000000 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=4 | DataOutVld=1 | RA=0 | CA=0 | cs_n=0
#                   55 | rst_n=1 | Addr=0000 | cmd_n=1 | RDnWR=0 | DataIn=00000000 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=1 | RA=0 | CA=0 | cs_n=0
#                   65 | rst_n=1 | Addr=0000 | cmd_n=1 | RDnWR=0 | DataIn=00000000 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=4 | DataOutVld=1 | RA=0 | CA=0 | cs_n=0
#                   75 | rst_n=1 | Addr=0000 | cmd_n=1 | RDnWR=0 | DataIn=00000000 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=1 | RA=0 | CA=0 | cs_n=0


# [WRITE] Addr: 1001, Data: a5a5a5a5
#                  245 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=0 | DataIn=a5a5a5a5 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=1 | DataOutVld=1 | RA=0 | CA=0 | cs_n=0
#                  255 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=0 | DataIn=a5a5a5a5 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  265 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=0 | DataIn=a5a5a5a5 | DQ=a5a5a5a5 | DataOut=00000000 | Cmd=3 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  275 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=0 | DataIn=a5a5a5a5 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  325 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=0 | DataIn=a5a5a5a5 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=4 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  335 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=0 | DataIn=a5a5a5a5 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  345 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=0 | DataIn=a5a5a5a5 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=4 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  355 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=0 | DataIn=a5a5a5a5 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0                425 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=0 | DataIn=a5a5a5a5 | DQ=zzzzzzzz | DataOut=00000000 | Cmd=4 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0

[WRITE] Addr: 2000, Data: deadbeef
#                  565 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=0 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=00000000 | Cmd=1 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  575 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=0 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=1 | RA=10 | CA=0 | cs_n=0
#                  635 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=0 | DataIn=deadbeef | DQ=deadbeef | DataOut=00000000 | Cmd=3 | DataOutVld=1 | RA=10 | CA=0 | cs_n=0
#                  645 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=0 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=00000000 | Cmd=0 | DataOutVld=1 | RA=10 | CA=0 | cs_n=0

# [READ] Addr: 1001, DataOut: 00000000, Valid: 1
#                  945 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=00000000 | Cmd=2 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  955 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=a5a5a5a5 | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  985 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=a5a5a5a5 | Cmd=2 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                  995 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=a5a5a5a5 | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0

# [READ] Addr: 2000, DataOut: deadbeef, Valid: 1
#                 1345 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=4 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                 1355 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                 1365 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=4 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                 1375 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0

# [READ] Addr: 1001, DataOut: deadbeef, Valid: 1
#                 2455 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                 2465 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=4 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                 2475 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                 2485 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=4 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                 2495 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=0 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0
#                 2505 | rst_n=1 | Addr=1001 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=deadbeef | Cmd=4 | DataOutVld=1 | RA=1 | CA=1 | cs_n=0


[READ] Addr: 2000, DataOut: 5a5a5a5b, Valid: 1
#                 3405 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=5a5a5a5b | Cmd=0 | DataOutVld=1 | RA=10 | CA=0 | cs_n=0
#                 3415 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=5a5a5a5b | Cmd=4 | DataOutVld=1 | RA=10 | CA=0 | cs_n=0
#                 3425 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=5a5a5a5b | Cmd=0 | DataOutVld=1 | RA=10 | CA=0 | cs_n=0
#                 3435 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=5a5a5a5b | Cmd=4 | DataOutVld=1 | RA=10 | CA=0 | cs_n=0
#                 3445 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=5a5a5a5b | Cmd=0 | DataOutVld=1 | RA=10 | CA=0 | cs_n=0
#                 3455 | rst_n=1 | Addr=2000 | cmd_n=1 | RDnWR=1 | DataIn=deadbeef | DQ=zzzzzzzz | DataOut=5a5a5a5b | Cmd=4 | DataOutVld=1 | RA=10 | CA=0 | cs_n=0