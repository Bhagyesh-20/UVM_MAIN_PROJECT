`include "interface.sv"
package pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    `include "transaction.sv"
    `include "rd_sequence.sv"
    `include "rst_sequence.sv"
    `include "wr_invld_sequence.sv"
    `include "randomize_sequence.sv"
    `include "wr_sequence.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "scoreboard.sv"
    `include "agent.sv"
    `include "env.sv"
    `include "test.sv"
endpackage
